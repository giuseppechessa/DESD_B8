library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity VolumeController.vhd is
	generic (
		NBITSNORMAL : INTEGER := 6
	);
	Port ( 
		aclk 			: in  STD_LOGIC;
		aresetn			: in  STD_LOGIC;

	);
end VolumeController.vhd;

architecture Behavioral of LED_Unpacker is


	
begin
    
     

end Behavioral;